`ifndef UVM_EXT_MONITOR_SV
	`define UVM_EXT_MONITOR_SV
	class uvm_ext_monitor#(type VIRTUAL_INTF=int,type ITEM_MON=uvm_sequence_item) extends uvm_monitor implements uvm_ext_reset_handler;
		
		uvm_ext_agent_config#(VIRTUAL_INTF) agent_config;
		
		protected process process_collect_transactions;

		uvm_analysis_port#(ITEM_MON) output_port; 

		`uvm_component_param_utils(uvm_ext_monitor#(VIRTUAL_INTF,ITEM_MON))

		function new(string name="",uvm_component parent);
			super.new(name,parent);
			output_port=new("output_port",this);
		endfunction : new

		virtual task wait_reset_end();
			agent_config.wait_reset_end();
		endtask : wait_reset_end
		
		virtual task run_phase(uvm_phase phase);
			forever begin
        		fork
          			begin
            			wait_reset_end();
            			collect_transactions();
            			disable fork;
          			end
        		join
      		end
		endtask : run_phase
     	
            

		protected virtual task collect_transactions();
			fork
				begin
					process_collect_transactions=process::self();
					begin
						forever begin
							collect_transaction();
						end
					end
				end	

			join		
		endtask : collect_transactions

		protected virtual task collect_transaction();
			`uvm_fatal("ALGORITHM_ISSUE","one must implement collect_transaction task()")
		endtask : collect_transaction

		virtual function void handle_reset(uvm_phase phase);
			if (process_collect_transactions!=null) begin
				process_collect_transactions.kill();
				process_collect_transactions=null;
			end
        endfunction

	endclass : uvm_ext_monitor
`endif